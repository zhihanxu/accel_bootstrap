module bank3_uram #(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 21
) (
    input clk,
    input [ADDR_WIDTH-1:0] addr,
    input [DATA_WIDTH-1:0] data_in,
    output reg [DATA_WIDTH-1:0] data_out,
    input we
);
    // Declare the URAM memory array
    (* ram_style = "ultra" *) reg [DATA_WIDTH-1:0] ram [0:(1<<ADDR_WIDTH)-1];

    always @(posedge clk) begin
        if (we) begin
            ram[addr] <= data_in;
        end
        data_out <= ram[addr];
    end
endmodule

module bank4_uram #(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 22
) (
    input clk,
    input [ADDR_WIDTH-1:0] addr,
    input [DATA_WIDTH-1:0] data_in,
    output reg [DATA_WIDTH-1:0] data_out,
    input we
);
    // Declare the URAM memory array
    (* ram_style = "ultra" *) reg [DATA_WIDTH-1:0] ram [0:(1<<ADDR_WIDTH)-1];

    always @(posedge clk) begin
        if (we) begin
            ram[addr] <= data_in;
        end
        data_out <= ram[addr];
    end
endmodule